module or_gate(a, b, out); //module is a keyword whereas or_gate is an identifier or name
input a,b;//input is a keyword
output out;//output is a keyword
or or1(out,a,b);
endmodule //or_gate